module proc(Data, Reset, w, Clock, F, Rx, Ry, Done, BusWires);
	input [7:0] Data;
	input Reset, w, Clock;
	input [1:0] F, Rx, Ry;
	output reg [7:0] BusWires;
	output reg Done;
	reg [7:0] Sum;
	reg [0:3] Rin, Rout;
	reg Extern, Ain, Gin, Gout, AddSub;
	wire [1:0] Count, I;
	wire [0:3] Xreg, Y;
	wire [7:0] R0, R1, R2, R3, A, G;
	wire [1:6] Func, FuncReg, Sel;
	
	wire Clear = Reset | Done | (~w & ~Count[1] & ~Count[0]);
	upcount counter (Clear, Clock, Count);
	assign Func = {F, Rx, Ry};
	wire FRin = w & ~Count[1] & ~Count[0];
	regn functionreg (Func, FRin, Clock, FuncReg);
		defparam functionreg.n = 6;
	assign I = FuncReg[1:2];
	dec2to4 decX (FuncReg[3:4], 1'b1, Xreg);
	dec2to4 decY (FuncReg[5:6], 1'b1, Y);

	always @(Count, I, Xreg , Y)
	begin
		Extern = 1'b0;  Done = 1'b0;  Ain = 1'b0;  Gin = 1'b0;
		Gout = 1'b0;  AddSub = 1'b0;  Rin = 4'b0;  Rout = 4'b0;
		case (Count)
			2'b00:	; // no signals asserted in time step T0
			2'b01:   // define signals in time step T1
						case (I)
							2'b00:	begin  //Load
											Extern = 1'b1;  Rin = Xreg;  Done = 1'b1;
										end
							2'b01:	begin  //Move
											Rout = Y; Rin = Xreg;  Done = 1'b1;
										end
							default: begin  //Add, Sub 
											Rout = Xreg; Ain = 1'b1;					            			 
					 					end		  
						endcase
         2'b10:	//define signals in time step T2
						case (I)
		           		2'b10: 	begin  //Add						           						
											Rout = Y; Gin = 1'b1;
							 			end
		              	2'b11: 	begin  //Sub		
			          					Rout = Y;  AddSub = 1'b1;  Gin = 1'b1;
										end
		    				default: ; //Add, Sub
						endcase
			2'b11: 
						case (I)
		    				2'b10, 2'b11:  begin
			           							Gout = 1'b1; Rin = Xreg; Done = 1'b1;
			      							end
		    				default: ; //Add, Sub
						endcase
	  	endcase
	end

	regn reg_0 (BusWires, Rin[0], Clock, R0);
	regn reg_1 (BusWires, Rin[1], Clock, R1);
	regn reg_2 (BusWires, Rin[2], Clock, R2);
	regn reg_3 (BusWires, Rin[3], Clock, R3);
	regn reg_A (BusWires, Ain, Clock, A);

	//alu
	always @(AddSub, A, BusWires)
	begin
	  	if (!AddSub)
		   Sum = A + BusWires;
    	else	
        	Sum = A - BusWires;
	end

	regn reg_G (Sum, Gin, Clock, G);
	assign Sel = {Rout, Gout, Extern};

	always @(Sel, R0,  R1, R2, R3, G, Data)
	begin
   	if (Sel == 6'b100000)
 			BusWires = R0;
  		else if (Sel == 6'b010000)
  			BusWires = R1;
  		else if (Sel == 6'b001000)
  			BusWires = R2;
  		else if (Sel == 6'b000100)
  			BusWires = R3;
  	 	else if (Sel == 6'b000010)
  			BusWires = G;
  		else BusWires = Data;
	end

endmodule
	

